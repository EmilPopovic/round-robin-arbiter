`timescale 1ns/1ps

module tb_round_robin_arbiter();

logic clk = 0;
logic rstn = 0;

endmodule
